library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.core_pack.all;
use work.fetch_pkg.all;

entity fetch_tb is
end fetch_tb;

architecture rtl of fetch_tb is
begin

end architecture rtl;