library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.core_pack.all;
use work.op_pack.all;

entity fwd is
	--port (
		-- define input and output ports as needed
--);
	
end fwd;

architecture rtl of fwd is

begin  -- rtl

end rtl;
