entity exec_tb is
end entity;

architecture rtl of exec_tb is
begin
end architecture;