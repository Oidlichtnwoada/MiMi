library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.core_pack.all;
use work.op_pack.all;

package decode_pkg is

    component decode is 
        port (
            clk, reset : in  std_logic;
            stall      : in  std_logic;
            flush      : in  std_logic;
            pc_in      : in  std_logic_vector(PC_WIDTH-1 downto 0);
            instr	   : in  std_logic_vector(INSTR_WIDTH-1 downto 0);
            wraddr     : in  std_logic_vector(REG_BITS-1 downto 0);
            wrdata     : in  std_logic_vector(DATA_WIDTH-1 downto 0);
            regwrite   : in  std_logic;
            pc_out     : out std_logic_vector(PC_WIDTH-1 downto 0);
            exec_op    : out exec_op_type;
            cop0_op    : out cop0_op_type;
            jmp_op     : out jmp_op_type;
            mem_op     : out mem_op_type;
            wb_op      : out wb_op_type;
            exc_dec    : out std_logic
        );
    end component;

end package;