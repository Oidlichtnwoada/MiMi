library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.core_pack.all;

entity regfile_tb is 
end regfile_tb;

architecture rtl of regfile_tb is 
begin
end rtl;