entity jmpu_tb is
end entity;

architecture rtl of jmpu_tb is
begin
end architecture;