library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.core_pack.all;

package fetch_pkg is

    component fetch is 
        port (
            clk, reset : in	 std_logic;
            stall      : in  std_logic;
            pcsrc	   : in	 std_logic;
            pc_in	   : in	 std_logic_vector(PC_WIDTH-1 downto 0);
            pc_out	   : out std_logic_vector(PC_WIDTH-1 downto 0);
            instr	   : out std_logic_vector(INSTR_WIDTH-1 downto 0)
        );
    end component;

end package;